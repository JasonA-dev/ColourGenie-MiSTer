//-------------------------------------------------------------------------------------------------
module clock
//-------------------------------------------------------------------------------------------------
(
	input  wire i, // 50.0000 MHz
	output wire o  // 35.4166 MHz (should be 35.4688 MHz, 17.7344*2)
);
//-------------------------------------------------------------------------------------------------

IBUFG IBufg(.I(i), .O(ci));

PLL_BASE #
(
	.CLKIN_PERIOD      (20.000),
	.CLKFBOUT_MULT     (17    ),
	.DIVCLK_DIVIDE     ( 1    ),
	.CLKOUT0_DIVIDE    (24    )
)
Pll
(
	.RST               (1'b0),
	.CLKFBIN           (fb),
	.CLKFBOUT          (fb),
	.CLKIN             (ci),
	.CLKOUT0           (co),
	.CLKOUT1           (),
	.CLKOUT2           (),
	.CLKOUT3           (),
	.CLKOUT4           (),
	.CLKOUT5           (),
	.LOCKED            ()
);

BUFG Bufg17(.I(co), .O(o));

//-------------------------------------------------------------------------------------------------
endmodule
//-------------------------------------------------------------------------------------------------
